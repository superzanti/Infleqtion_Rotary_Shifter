LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY fpga_top IS

END ENTITY fpga_top;

ARCHITECTURE rtl OF fpga_top IS

BEGIN

END ARCHITECTURE rtl;